package yapp_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "yapp_packet.sv"
    `include "router_tb.sv"
    `include "router_test_lib.sv"

endpackage : yapp_pkg